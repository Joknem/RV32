`include "../core/defines.v"

module gpio (
    input wire clk,
    input wire rst,
);
endmodule