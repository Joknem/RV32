`include "../core/defines.v"

module bus(
    input wire clk,
    input wire rst,
    input wire slave_
);
endmodule